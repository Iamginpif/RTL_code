package fa_package;
    `include "full_adder.sv"
    `include "add_subtract.sv"
endpackage

